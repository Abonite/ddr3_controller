library IEEE;

use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity write_levleing is
    port(
        clk : in std_logic;
        
        start_write_leveling : in std_logic
    );
end entity write_levleing;

architecture Behavioral of write_levleing is
    
begin
    
end architecture Behavioral;

